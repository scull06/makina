module alu16 (
    input wire [15:0] A,
    input wire [15:0] B,
    input wire [7:0] ALUop,
    output wire [15:0] Result
);
    
endmodule



module adder16 (
    input wire  [15:0] A,
    input wire  [15:0] B,
    output wire [15:0] Result
);

 
    
endmodule